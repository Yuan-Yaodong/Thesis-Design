module UCAC3(
    input x1,
    input x2,
    input x3,
    input x4,
    output sum
);

    assign sum = x2 | x4;

endmodule
