
module AHA(
    input x1,
    input x2,
    output sum
);

    assign sum = x1 | x2;

endmodule

